module ADDER_FOUR(
input [31:0] ADDER_FOUR_IN,
output [31:0] ADDER_FOUR_OUT
);

assign  ADDER_FOUR_OUT = ADDER_FOUR_IN + 4;


endmodule